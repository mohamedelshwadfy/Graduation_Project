/* Module: CarryLookAhead4Bit
   Description: 4-bit Carry Look-Ahead Adder
   Inputs: a, b - 4-bit input lines; cin - Carry input
   Outputs: sum - 4-bit sum; cout - Carry output
*/
module CarryLookAhead4Bit ( 
    input  [3:0]  a,
    input  [3:0]  b,
    input         cin,
    output [3:0]  sum,
    output        cout
);
    wire   [3:0]  p;
    wire   [3:0]  g;
    wire   [3:0]  c;

    assign p = a ^ b;      // propagate
    assign g = a & b;      // generate
    assign c[0] = cin;
    assign c[1] = g[0] | (p[0] & c[0]);
    assign c[2] = g[1] | (p[1] & g[0]) | (p[1] & p[0] & c[0]);
    assign c[3] = g[2] | (p[2] & g[1]) | (p[2] & p[1] & g[0]) | (p[2] & p[1] & p[0] & c[0]);
    assign cout = g[3] | (p[3] & g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0]) | (p[3] & p[2] & p[1] & p[0] & c[0]);
    assign sum = p ^ c;

endmodule

